`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:44:52 06/01/2016 
// Design Name: 
// Module Name:    denormalization_module 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module denormalization_module(
    input [39:0] operand,
    input type_shift,
    output [31:0] denorm_operand
    );


endmodule
